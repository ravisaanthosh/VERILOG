module rc(input clk,rs,output reg [3:0]q);
always @(posedge clk)begin
if(rs==0)
q<=4'b1110;
else begin
q[3]<=q[0];
q[2]<=q[3];
q[1]<=q[2];
q[0]<=q[1];
end
end
endmodule

