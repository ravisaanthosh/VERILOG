

//D RAM HAVE A PERIODIC REFRESH TO PTORECT A DATA HERE WE CAN'T ADD A PERIODIC REFRESH IN CODING ITS A HARDWARE COMPONENTS AND SAME AS A S RAM SINGLE PORT ,, D RAM ONLY AVIALABE IN SINGLE PORT ONLY 
module Dram(input clk,rs,wr,input[3:0]din,input[2:0]add,output reg[3:0]dout);
reg[7:0] ram[3:0];   //7:0 represents in adderess 3:0 represents in data
always@(posedge clk)begin
//reset purpose
if(rs==1)
dout<=4'b0000;
//write purpose
else if(wr==1)
ram[add]<=din;
//read purpose
else if(wr==0)
dout<=ram[add];
end
endmodule
