module epg(input a,b,c,output p);
assign p=(a^b^c);
endmodule
